CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 146 195 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5476 0 0
2
5.89884e-315 0
0
9 CC 7-Seg~
183 998 130 0 18 19
10 11 10 9 8 7 6 5 18 19
0 0 0 0 0 0 0 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3936 0 0
2
5.89884e-315 5.26354e-315
0
9 2-In AND~
219 539 46 0 3 22
0 15 3 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5770 0 0
2
5.89884e-315 5.30499e-315
0
9 2-In AND~
219 400 36 0 3 22
0 4 13 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7884 0 0
2
5.89884e-315 5.32571e-315
0
6 74112~
219 604 225 0 7 32
0 17 14 16 14 17 20 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3690 0 0
2
5.89884e-315 5.34643e-315
0
6 74112~
219 504 226 0 7 32
0 17 15 16 15 17 21 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3611 0 0
2
5.89884e-315 5.3568e-315
0
6 74112~
219 395 231 0 7 32
0 17 4 16 4 17 22 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7912 0 0
2
5.89884e-315 5.36716e-315
0
6 74112~
219 289 231 0 7 32
0 17 2 16 2 17 23 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6416 0 0
2
5.89884e-315 5.37752e-315
0
6 74LS48
188 845 204 0 14 29
0 12 3 13 4 24 25 5 6 7
8 9 10 11 26
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7278 0 0
2
5.89884e-315 5.38788e-315
0
2 +V
167 145 123 0 1 3
0 17
0
0 0 54256 0
2 5V
-6 -22 8 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6804 0 0
2
5.89884e-315 5.39306e-315
0
7 Pulser~
4 145 312 0 10 12
0 27 28 16 29 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9568 0 0
2
5.89884e-315 5.39824e-315
0
35
4 0 2 0 0 4096 0 8 0 0 2 3
265 213
172 213
172 195
1 2 2 0 0 4224 0 1 8 0 0 2
158 195
265 195
2 0 3 0 0 12416 0 9 0 0 17 4
813 177
784 177
784 151
512 151
0 2 4 0 0 4096 0 0 7 26 0 2
343 195
371 195
7 7 5 0 0 4224 0 9 2 0 0 3
877 168
1013 168
1013 166
8 6 6 0 0 4224 0 9 2 0 0 3
877 177
1007 177
1007 166
9 5 7 0 0 4224 0 9 2 0 0 3
877 186
1001 186
1001 166
10 4 8 0 0 4224 0 9 2 0 0 3
877 195
995 195
995 166
11 3 9 0 0 4224 0 9 2 0 0 3
877 204
989 204
989 166
4 7 4 0 0 8320 0 9 8 0 0 5
813 195
813 288
327 288
327 195
313 195
12 2 10 0 0 4224 0 9 2 0 0 3
877 213
983 213
983 166
13 1 11 0 0 4224 0 9 2 0 0 3
877 222
977 222
977 166
7 1 12 0 0 4224 0 5 9 0 0 4
628 189
803 189
803 168
813 168
0 3 13 0 0 4224 0 0 9 21 0 4
433 243
803 243
803 186
813 186
0 4 14 0 0 4224 0 0 5 16 0 3
566 95
566 207
580 207
3 2 14 0 0 0 0 3 5 0 0 5
560 46
560 95
566 95
566 189
580 189
2 7 3 0 0 0 0 3 6 0 0 6
515 55
512 55
512 159
539 159
539 190
528 190
0 4 15 0 0 4224 0 0 6 20 0 3
429 52
429 208
480 208
0 1 15 0 0 0 0 0 3 20 0 3
465 52
465 37
515 37
3 2 15 0 0 0 0 4 6 0 0 6
421 36
429 36
429 52
466 52
466 190
480 190
2 7 13 0 0 0 0 4 7 0 0 6
376 45
356 45
356 248
433 248
433 195
419 195
1 0 4 0 0 0 0 4 0 0 10 4
376 27
335 27
335 195
327 195
3 0 16 0 0 8192 0 5 0 0 24 4
574 198
570 198
570 302
470 302
3 0 16 0 0 12288 0 6 0 0 25 4
474 199
470 199
470 303
361 303
3 0 16 0 0 12416 0 7 0 0 27 4
365 204
361 204
361 304
251 304
0 4 4 0 0 0 0 0 7 22 0 4
335 195
343 195
343 213
371 213
3 3 16 0 0 128 0 11 8 0 0 6
169 303
251 303
251 304
251 304
251 204
259 204
5 0 17 0 0 8192 0 8 0 0 31 3
289 243
289 272
395 272
5 0 17 0 0 12288 0 5 0 0 32 5
604 237
604 272
668 272
668 134
602 134
5 0 17 0 0 0 0 6 0 0 29 3
504 238
504 272
604 272
5 0 17 0 0 0 0 7 0 0 30 3
395 243
395 272
504 272
0 1 17 0 0 0 0 0 5 33 0 3
504 134
604 134
604 162
0 1 17 0 0 0 0 0 6 34 0 3
395 134
504 134
504 163
1 0 17 0 0 0 0 7 0 0 35 3
395 168
395 134
289 134
1 1 17 0 0 4224 0 10 8 0 0 3
145 132
289 132
289 168
1
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 22
168 354 328 381
180 362 315 381
22 Hilot, Renalyn Bajenio
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
